--*****************************************************
--* Project ILECT
--* (c) copyright 2016
--* Company Magnetische Pruefanlagen GmbH
--* All rights reserved
--* Secrecy Level STRICTLY CONFIDENTIAL
--*****************************************************

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

library UNISIM;
use UNISIM.VComponents.all;

Library UNIMACRO;
use UNIMACRO.vcomponents.all;

entity packetRAM is
      -- NB! Memory Size is 36Kbits
      generic (
         g_port1_dat_width : natural := 32;
         g_port1_adr_width : natural := 9;
         g_port2_dat_width : natural := 32;
         g_port2_adr_width : natural := 9
         
         );
      port (
         i_clk1 : in  std_logic;
         i_rst1 : in  std_logic;
         i_wre1 : in  std_logic;
         i_dat1 : in  std_logic_vector(g_port1_dat_width - 1 downto 0);
         i_adr1 : in  std_logic_vector(g_port1_adr_width - 1 downto 0);

         i_clk2 : in  std_logic;
         i_rst2 : in  std_logic;
         i_rde2 : in  std_logic;
         o_dat2 : out std_logic_vector(g_port2_dat_width - 1 downto 0);
         i_adr2 : in  std_logic_vector(g_port2_adr_width - 1 downto 0)
      );

end packetRAM;

architecture Behavioral of packetRAM is
      constant s_ones   : std_logic_vector(31 downto 0) := X"FFFF_FFFF";
      constant s_zeros  : std_logic_vector(31 downto 0) := X"0000_0000";
begin   
   -- BRAM_TDP_MACRO: True Dual Port RAM
   --                 Artix-7
   -- Xilinx HDL Language Template, version 2016.2

   -- Note -  This Unimacro model assumes the port directions to be "downto". 
   --         Simulation of this model with "to" in the port directions could lead to erroneous results.

   --------------------------------------------------------------------------
   -- DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width --
   -- ===============|===========|===========|===============|=============--
   --     19-36      |  "36Kb"   |    1024   |    10-bit     |    4-bit    --
   --     10-18      |  "36Kb"   |    2048   |    11-bit     |    2-bit    --
   --     10-18      |  "18Kb"   |    1024   |    10-bit     |    2-bit    --
   --      5-9       |  "36Kb"   |    4096   |    12-bit     |    1-bit    --
   --      5-9       |  "18Kb"   |    2048   |    11-bit     |    1-bit    --
   --      3-4       |  "36Kb"   |    8192   |    13-bit     |    1-bit    --
   --      3-4       |  "18Kb"   |    4096   |    12-bit     |    1-bit    --
   --        2       |  "36Kb"   |   16384   |    14-bit     |    1-bit    --
   --        2       |  "18Kb"   |    8192   |    13-bit     |    1-bit    --
   --        1       |  "36Kb"   |   32768   |    15-bit     |    1-bit    --
   --        1       |  "18Kb"   |   16384   |    14-bit     |    1-bit    --
   --------------------------------------------------------------------------
   
   BRAM_TDP_MACRO_inst : BRAM_TDP_MACRO
   generic map (
      BRAM_SIZE         => "36Kb", -- Target BRAM, "18Kb" or "36Kb" 
      DEVICE            => "7SERIES", -- Target Device: "VIRTEX5", "VIRTEX6", "7SERIES", "SPARTAN6" 
      DOA_REG           => 0, -- Optional port A output register (0 or 1)
      DOB_REG           => 0, -- Optional port B output register (0 or 1)
      INIT_A            => X"000000000", -- Initial values on A output port
      INIT_B            => X"000000000", -- Initial values on B output port
      INIT_FILE         => "NONE",
      READ_WIDTH_A      => g_port1_dat_width,   -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
      READ_WIDTH_B      => g_port2_dat_width,   -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
      SIM_COLLISION_CHECK => "ALL", -- Collision check enable "ALL", "WARNING_ONLY", 
                                    -- "GENERATE_X_ONLY" or "NONE" 
      SRVAL_A           => X"000000000",   -- Set/Reset value for A port output
      SRVAL_B           => X"000000000",   -- Set/Reset value for B port output
      WRITE_MODE_A      => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE" 
      WRITE_MODE_B      => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE" 
      WRITE_WIDTH_A     => g_port1_dat_width, -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
      WRITE_WIDTH_B     => g_port2_dat_width, -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
      -- The following INIT_xx declarations specify the initial contents of the RAM
      INIT_00           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F           => X"0000000000000000000000000000000000000000000000000000000000000000",
      
      -- The next set of INIT_xx are valid when configured as 36Kb
      INIT_40           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_41           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_42           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_43           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_44           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_45           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_46           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_47           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_48           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_49           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4A           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4B           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4C           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4D           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4E           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4F           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_50           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_51           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_52           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_53           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_54           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_55           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_56           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_57           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_58           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_59           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5A           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5B           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5C           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5D           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5E           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5F           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_60           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_61           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_62           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_63           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_64           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_65           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_66           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_67           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_68           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_69           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6A           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6B           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6C           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6D           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6E           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6F           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_70           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_71           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_72           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_73           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_74           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_75           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_76           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_77           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_78           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_79           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7A           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7B           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7C           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7D           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7E           => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7F           => X"0000000000000000000000000000000000000000000000000000000000000000",
      
      -- The next set of INITP_xx are for the parity bits
      INITP_00          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07          => X"0000000000000000000000000000000000000000000000000000000000000000",
      
      -- The next set of INIT_xx are valid when configured as 36Kb
      INITP_08          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_09          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0A          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0B          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0C          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0D          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0E          => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0F          => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA               => open,             -- Output port-A data, width defined by READ_WIDTH_A parameter
      DOB               => o_dat2,           -- Output port-B data, width defined by READ_WIDTH_B parameter
      ADDRA             => i_adr1,           -- Input port-A address, width defined by Port A depth
      ADDRB             => i_adr2,           -- Input port-B address, width defined by Port B depth
      CLKA              => i_clk1,           -- 1-bit input port-A clock
      CLKB              => i_clk2,           -- 1-bit input port-B clock
      DIA               => i_dat1,           -- Input port-A data, width defined by WRITE_WIDTH_A parameter
      DIB               => (others => '0'),  -- Input port-B data, width defined by WRITE_WIDTH_B parameter
      ENA               => i_wre1,           -- 1-bit input port-A enable
      ENB               => i_rde2,           -- 1-bit input port-B enable
      REGCEA            => '1',              -- 1-bit input port-A output register enable
      REGCEB            => '1',              -- 1-bit input port-B output register enable
      RSTA              => i_rst1,              -- 1-bit input port-A reset
      RSTB              => i_rst2,              -- 1-bit input port-B reset
      WEA               => s_ones(g_port1_dat_width / 8  - 1 downto 0),  -- Input port-A write enable, width defined by Port A depth
      WEB               => s_zeros(g_port2_dat_width / 8  - 1 downto 0)   -- Input port-B write enable, width defined by Port B depth
   );
   
end Behavioral;
